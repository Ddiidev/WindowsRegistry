module winreg

pub enum Reserved as u32 {
	rrf_rt_reg_dword = 0x00000010
}
