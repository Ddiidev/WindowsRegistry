module winreg

pub struct InfoValues {
pub mut:
	name string
	typ  DwType
}
